module tb;
    reg [63:0] x;             
    integer i;
    reg [63:0] pattern [0:31]; 
    initial begin
       
        pattern[0]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        pattern[1]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        pattern[2]  = 64'b0000000000000000000000000000000000000000000000000000000000000000; 
        pattern[3]  = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        pattern[4]  = 64'b0000000000000000000000100100000000000000000000000000000000001111;
        pattern[5]  = 64'b0000000000000000000001110100000000000000000000000000000000001111;
        pattern[6]  = 64'b0000000000000000000011111100000000000000000000011111110000001111; 
        pattern[7]  = 64'b0000000000000000000001110100001111111111111000100000001000001111;
        pattern[8]  = 64'b0001111111111110000000100100010000000000000100100000000100001111;
        pattern[9]  = 64'b0010000000000001000000000100100000000000000010010000000100001111;
        pattern[10]  = 64'b0100000000000010000011111101000000000000000001010000000010001111; 
        pattern[11]  = 64'b0010000000000100000100000010000000000000000000110000000010001111;
        pattern[12]  = 64'b0001000000001000001000000010000000000000000000010000000010001111;
        pattern[13]  = 64'b0000111111111000010000000000000000000000000000010000000010001111;
        pattern[14]  = 64'b0001000000000100100000000000000000000000000000010000000010001111;
        pattern[15]  = 64'b0011000000000010100000000000001100000000000000010000000001111111; 
        pattern[16]  = 64'b0111000100000001000000000000000010000000000000010000000000111111;
        pattern[17]  = 64'b1111000000000000111111111111111100000000000000010000000000011111;
        pattern[18]  = 64'b0111000100000001000000000000000000000000000000010000000111101111;
        pattern[19]  = 64'b0011000000000010100000000000000000000000000000010000001000001111; 
        pattern[20]  = 64'b0001000000000100010000000000000000000000000000010000000100001111;
        pattern[21]  = 64'b0000111111111000001000000010000000000000000000010000000010001111;
        pattern[22]  = 64'b0001000000001000000100000010000000000000000000110000000010001111;
        pattern[23]  = 64'b0010000000000100000001111101000000000000000001010000000010001111; 
        pattern[24]  = 64'b0100000000000010000000000010100000000000000010010000000010001111;
        pattern[25]  = 64'b0100000000000001000000111110010000000000000100100000000010001111;
        pattern[26]  = 64'b0011111111111110000000111110001111111111111001000000000100001111;
        pattern[27]  = 64'b0000000000000000000000000010000000000000000000100000000100001111; 
        pattern[28]  = 64'b0000000000000000000000000000000000000000000000100000001000001111;
        pattern[29]  = 64'b0000000000000000000000000000000000000000000000011111110000001111;
        pattern[30]  = 64'b0000000000000000000000000000000000000000000000000000000000001111;
        pattern[31]  = 64'b0000000000000000000000000000000000000000000000000000000100001111; 
        
 
 
        for (i = 0; i < 45; i = i + 1) begin
            x = pattern[i];
            #10; // 10ns per step
        end
        $finish;
    end
endmodule
