// Code your testbench here
// or browse Examples
module tb ;
  reg [0:10]a;
  initial 
    begin
      $dumpfile("dump.vcd"); $dumpvars;
      a=11'b00000000000;#5;
      a=11'b11111111111;#5;
      a=11'b00000100000;#5;
      a=11'b00000100000;#5;
      a=11'b11111111111;#5;
      a=11'b00000000000;#5;
      a=11'b00011111111;#5;
      a=11'b01100010000;#5;
      a=11'b10000010000;#5;
      a=11'b01100010000;#5;
      a=11'b00011111111;#5;
      a=11'b00000000000;#5;
      a=11'b11111111111;#5;
      a=11'b10001000000;#5;
      a=11'b10001000000;#5;
      a=11'b01110000000;#5;
      a=11'b00000000000;#5;
      a=11'b11111111111;#5;
      a=11'b10001000000;#5;
      a=11'b10001000000;#5;
      a=11'b01110000000;#5;
      a=11'b00000000000;#5;
      a=11'b11000000100;#5;
      a=11'b00100000010;#5;
      a=11'b00010000001;#5;
      a=11'b11111111110;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b10000000000;#5;
      a=11'b10000000000;#5;
      a=11'b11111111111;#5;
      a=11'b10000000000;#5;      
      a=11'b10000000000;#5;
      a=11'b00000000000;#5;
      a=11'b11111111111;#5;
      a=11'b10000100001;#5;
      a=11'b10000100001;#5;      
      a=11'b10000000001;#5;
      a=11'b00000000000;#5;
      a=11'b00011111111;#5;
      a=11'b01100010000;#5;
      a=11'b10000010000;#5;
      a=11'b01100010000;#5;
      a=11'b00011111111;#5;
      a=11'b00000000000;#5;      
      a=11'b11111111111;#5;
      a=11'b10000000001;#5;
      a=11'b10000000001;#5;
      a=11'b10000000001;#5;
      a=11'b00000000000;#5;      
      a=11'b11111111111;#5;
      a=11'b00000100000;#5;
      a=11'b00000100000;#5;
      a=11'b11111111111;#5;
      a=11'b00000000000;#5;
      a=11'b11111111111;#5;
      a=11'b10000100001;#5;
      a=11'b10000100001;#5;      
      a=11'b10000000001;#5;
      a=11'b00000000000;#5;
      a=11'b11111111111;#5;
      a=11'b10001100000;#5;
      a=11'b10001010000;#5;
      a=11'b01110001111;#5;
      a=11'b00000000000;#5;      
      a=11'b11111100001;#5;
      a=11'b10000100001;#5;
      a=11'b10000100001;#5;
      a=11'b10000111111;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b11111111111;#5;
      a=11'b10000000001;#5;      
      a=11'b10000000001;#5;
      a=11'b01111111110;#5;
      a=11'b00000000000;#5;
      a=11'b00011111111;#5;
      a=11'b01100010000;#5;
      a=11'b10000010000;#5;
      a=11'b01100010000;#5;
      a=11'b00011111111;#5;
      a=11'b00000000000;#5;
      a=11'b11000000100;#5;
      a=11'b00100000010;#5;
      a=11'b00010000001;#5;
      a=11'b11111111110;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;      
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      a=11'b00000000000;#5;
      
    end
endmodule
